library verilog;
use verilog.vl_types.all;
entity system_hdmi_out_0_wrapper is
    port(
        PXL_CLK_X1      : in     vl_logic;
        PXL_CLK_X2      : in     vl_logic;
        PXL_CLK_X10     : in     vl_logic;
        PXL_PLL_LOCKED  : in     vl_logic;
        TMDS            : out    vl_logic_vector(3 downto 0);
        TMDSB           : out    vl_logic_vector(3 downto 0);
        S_AXI_ACLK      : in     vl_logic;
        S_AXI_ARESETN   : in     vl_logic;
        S_AXI_AWADDR    : in     vl_logic_vector(31 downto 0);
        S_AXI_AWVALID   : in     vl_logic;
        S_AXI_WDATA     : in     vl_logic_vector(31 downto 0);
        S_AXI_WSTRB     : in     vl_logic_vector(3 downto 0);
        S_AXI_WVALID    : in     vl_logic;
        S_AXI_BREADY    : in     vl_logic;
        S_AXI_ARADDR    : in     vl_logic_vector(31 downto 0);
        S_AXI_ARVALID   : in     vl_logic;
        S_AXI_RREADY    : in     vl_logic;
        S_AXI_ARREADY   : out    vl_logic;
        S_AXI_RDATA     : out    vl_logic_vector(31 downto 0);
        S_AXI_RRESP     : out    vl_logic_vector(1 downto 0);
        S_AXI_RVALID    : out    vl_logic;
        S_AXI_WREADY    : out    vl_logic;
        S_AXI_BRESP     : out    vl_logic_vector(1 downto 0);
        S_AXI_BVALID    : out    vl_logic;
        S_AXI_AWREADY   : out    vl_logic;
        m_axi_aclk      : in     vl_logic;
        m_axi_aresetn   : in     vl_logic;
        md_error        : out    vl_logic;
        m_axi_arready   : in     vl_logic;
        m_axi_arvalid   : out    vl_logic;
        m_axi_araddr    : out    vl_logic_vector(31 downto 0);
        m_axi_arlen     : out    vl_logic_vector(7 downto 0);
        m_axi_arsize    : out    vl_logic_vector(2 downto 0);
        m_axi_arburst   : out    vl_logic_vector(1 downto 0);
        m_axi_arprot    : out    vl_logic_vector(2 downto 0);
        m_axi_arcache   : out    vl_logic_vector(3 downto 0);
        m_axi_rready    : out    vl_logic;
        m_axi_rvalid    : in     vl_logic;
        m_axi_rdata     : in     vl_logic_vector(31 downto 0);
        m_axi_rresp     : in     vl_logic_vector(1 downto 0);
        m_axi_rlast     : in     vl_logic;
        m_axi_awready   : in     vl_logic;
        m_axi_awvalid   : out    vl_logic;
        m_axi_awaddr    : out    vl_logic_vector(31 downto 0);
        m_axi_awlen     : out    vl_logic_vector(7 downto 0);
        m_axi_awsize    : out    vl_logic_vector(2 downto 0);
        m_axi_awburst   : out    vl_logic_vector(1 downto 0);
        m_axi_awprot    : out    vl_logic_vector(2 downto 0);
        m_axi_awcache   : out    vl_logic_vector(3 downto 0);
        m_axi_wready    : in     vl_logic;
        m_axi_wvalid    : out    vl_logic;
        m_axi_wdata     : out    vl_logic_vector(31 downto 0);
        m_axi_wstrb     : out    vl_logic_vector(3 downto 0);
        m_axi_wlast     : out    vl_logic;
        m_axi_bready    : out    vl_logic;
        m_axi_bvalid    : in     vl_logic;
        m_axi_bresp     : in     vl_logic_vector(1 downto 0)
    );
end system_hdmi_out_0_wrapper;
